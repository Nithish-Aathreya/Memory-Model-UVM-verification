interface rintf(input bit clk);
  
  bit rst;
  bit [15:0] addr;
  bit wren;
  bit [7:0] wdata;
  bit [7:0]rdata;
  
  
  
  
  
  
endinterface
  
